`define DELAY 20
module ALU32_testbench(); 
reg [31:0] input1, input2;
reg [3:0] select;
reg carry_in;
wire carry_out_forAdd, carry_out_forSub;
wire [31:0] result;

ALU_32 test_ALU(result,carry_out_forAdd,carry_out_forSub,input1,input2,select,carry_in);

initial begin
input1 = 32'b11111111111111111111111111111111; input2 = 32'b00000000000000000000000000000000; select = 3'b000;
#`DELAY;
input1 = 32'b11111111111111111111111111111111; input2 = 32'b11111111111111111111111111111111; select = 3'b000;
#`DELAY;
input1 = 32'b01011010110101110110110101101011; input2 = 32'b00110000110101100100111101100001; select = 3'b000;
#`DELAY;
input1 = 32'b11111111111111111111111111111111; input2 = 32'b00000000000000000000000000000000; select = 3'b001;
#`DELAY;
input1 = 32'b00000000000000000000000000000000; input2 = 32'b00000000000000000000000000000000; select = 3'b001;
#`DELAY;
input1 = 32'b01011010110101110110110101101011; input2 = 32'b00110000110101100100111101100001; select = 3'b001;
#`DELAY;
input1 = 32'b11111111111111111111111111111111; input2 = 32'b11111111111111111111111111111111; select = 3'b010; carry_in = 1'b0;
#`DELAY;
input1 = 32'b11111111111111111111111111111111; input2 = 32'b00000000000000000000000000000000; select = 3'b010; carry_in = 1'b1;
#`DELAY;
input1 = 32'b00000000000000000000000000000000; input2 = 32'b00000000000000000000000000000000; select = 3'b010; carry_in = 1'b1;
#`DELAY;
input1 = 32'b10000010010101001100010000100010; input2 = 32'b00000010000001000011110000000001; select = 3'b011; 
#`DELAY;
input1 = 32'b10111100000000000010000001001001; input2 = 32'b01000010010000000000001000010001; select = 3'b011;
#`DELAY;
input1 = 32'b11001010101101111100011101010111; input2 = 32'b00101000000001110000000001111000; select = 3'b011; 
#`DELAY;
input1 = 32'b11111111111111111111111111111111; input2 = 32'b00000000000000000000000000000000; select = 3'b100; 
#`DELAY;
input1 = 32'b11111111111111111111111111111111; input2 = 32'b11111111111111111111111111111111; select = 3'b100; 
#`DELAY;
input1 = 32'b11111111111111111111111111100000; input2 = 32'b00000000000000000000000000011111; select = 3'b100;
#`DELAY;
input1 = 32'b10000000000000000000000100010000; input2 = 32'b00000000000000000000000000000011; select = 3'b101;
#`DELAY;
input1 = 32'b00000000000000000000100000000000; input2 = 32'b00000000000000000000000000001001; select = 3'b101;
#`DELAY;
input1 = 32'b10000000000000000000001100010000; input2 = 32'b00000000000000000000000000010101; select = 3'b101;
#`DELAY;
input1 = 32'b11111111111111111111111111111111; input2 = 32'b00000000000000000000000000000100; select = 3'b110; 
#`DELAY;
input1 = 32'b11111111111111000011111110110111; input2 = 32'b00000000000000000000000000001100; select = 3'b110; 
#`DELAY;
input1 = 32'b11111111111111111111111111111111; input2 = 32'b00000000000000000000000000011111; select = 3'b110; 
#`DELAY;
input1 = 32'b11000111111101111011101110111111; input2 = 32'b10001000000100010000010101010100; select = 3'b111; 
#`DELAY;
input1 = 32'b11001000100001000011101110110111; input2 = 32'b11000000110110101111010000001100; select = 3'b111; 
#`DELAY;
input1 = 32'b11110101111010000010011110111101; input2 = 32'b00111011010000011000001000011011; select = 3'b111; 
#`DELAY;
end
 
 
initial
begin

$monitor("time = %2d, input1 = %32b, input2 = %32b, select = %3b, result = %32b, carry_in = %1b, carry_out= %1b", $time, input1, input2, select, result, carry_in, carry_out_forAdd);

end
 
endmodule