`define DELAY 20
module LEFT_SHIFTER_testbench();
reg [31:0] input1, input2;
wire [31:0] result;

LEFT_SHIFTER f(result,input1,input2);
initial begin
input1 = 32'b00000000000000000000000000000011; input2 = 32'b00000000000000000000000000000001;
#`DELAY;
input1 = 32'b00000000000000000000000000000011; input2 = 32'b00000000000000000000000000000010;
#`DELAY;
input1 = 32'b00000000000000000000000000000011; input2 = 32'b00000000000000000000000000000011;
#`DELAY;
input1 = 32'b00000000000000000000000000000001; input2 = 32'b00000000000000000000000000011111;
#`DELAY;
input1 = 32'b00000000000000000000000000000001; input2 = 32'b00000000000000000000000000010000;
#`DELAY;
end 

initial
begin
$monitor("time = %2d, input1 = %32b, input2 = %32b,result = %32b", $time, input1, input2,result);
end

endmodule
